----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/14/2017 03:14:52 PM
-- Design Name: 
-- Module Name: inverter_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity inverter_tb is
--  Port ( );
end inverter_tb;

architecture Behavioral of inverter_tb is
--signal input, output: std_logic_vector(1 downto 0);
--begin
--some: entity work.inverter port map(sw=>input,led=>output);
----some_2: entity work.inverter port map(b=>input,a=>output);
--stimulus: process
--begin
--input<="01";
--wait for 100 ns;
--input<="10";
--wait for 100 ns;

--end process;

--some: entity work.inverter port map(a=>input,b=>output);

end Behavioral;
